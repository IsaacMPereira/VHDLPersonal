library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity judges_ex5 is
    Port ( a, b, c, d : in STD_LOGIC;
           m, u, c : out STD_LOGIC);
end judges_ex5;

architecture Behavioral of judges_ex5 is

begin
    
end Behavioral;
